library ieee;
   use ieee.std_logic_1164.all;


package wbfbd is

   type t_slv_vector is array (natural range <>) of std_logic_vector;

   type t_integer_vector is array (natural range <>) of integer;

   -- FBDL main package and main bus constants.
{Constants}
end package;
